module dFF #(parameter n = 32) (
  input  logic          clk,
  input  logic          reset,
  input  logic [n-1:0]  d,
  output logic [n-1:0]  q
);

always_ff @(posedge clk) begin
  if (reset)  q <= 0;
  else        q <= d;
end

endmodule